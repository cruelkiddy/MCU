library verilog;
use verilog.vl_types.all;
entity MCU2_vlg_vec_tst is
end MCU2_vlg_vec_tst;
